// Author: Shane Nelson
// Project: OoO CPU
// File: IF to Issue pipeline register
// Stage: Fetch -> Issue

module pipeline_reg (
    input  pipe_in_t d,
    input  logic reset, clk, queue_full,
    output pipe_in_t q
);
    pipe_in_t q_reg;

    assign q = q_reg;

    always_ff @(posedge clk) begin
        if (reset) begin  // flush reg on reset or flush
            q_reg.instruction <= 32'b0;
            q_reg.pc <= 32'b0;
            q_reg.prediction  <= 1'b0;
        end
        else if (!queue_full) begin  // if issue queue can accept new data, update
            q_reg <= d;
        end
    end
endmodule